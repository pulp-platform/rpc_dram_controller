// rpc top module for fpga synthesis

module rpc_xilinx (

    // clock and reset
    input  wire             clkp_i,
    input  wire             clkn_i,
    input  wire             rst_ni,

    // axi slave interface
    input  [ 5:0]           axi_aw_id_i,
    input  [ 39:0]          axi_aw_addr_i,
    input  [ 7:0]           axi_aw_len_i,
    input  [ 2:0]           axi_aw_size_i,
    input  [ 1:0]           axi_aw_burst_i,
    input                   axi_aw_lock_i,
    input  [ 3:0]           axi_aw_cache_i,
    input  [ 2:0]           axi_aw_prot_i,
    input  [ 3:0]           axi_aw_qos_i,
    input  [ 3:0]           axi_aw_region_i,
    input  [ 5:0]           axi_aw_atop_i,
    input                   axi_aw_user_i,
    input                   axi_aw_valid_i,
    output                  axi_aw_ready_o,
    input  [ 63:0]          axi_w_data_i,
    input  [ 7:0]           axi_w_strb_i,
    input                   axi_w_last_i,
    input                   axi_w_user_i,
    input                   axi_w_valid_i,
    output                  axi_w_ready_o,
    output [ 5:0]           axi_b_id_o,
    output [ 1:0]           axi_b_resp_o,
    output                  axi_b_user_o,
    output                  axi_b_valid_o,
    input                   axi_b_ready_i,
    input  [ 5:0]           axi_ar_id_i,
    input  [ 39:0]          axi_ar_addr_i,
    input  [ 7:0]           axi_ar_len_i,
    input  [ 2:0]           axi_ar_size_i,
    input  [ 1:0]           axi_ar_burst_i,
    input                   axi_ar_lock_i,
    input  [ 3:0]           axi_ar_cache_i,
    input  [ 2:0]           axi_ar_prot_i,
    input  [ 3:0]           axi_ar_qos_i,
    input  [ 3:0]           axi_ar_region_i,
    input  [ 0:0]           axi_ar_user_i,
    input                   axi_ar_valid_i,
    output                  axi_ar_ready_o,
    output [ 5:0]           axi_r_id_o,
    output [ 63:0]          axi_r_data_o,
    output [ 1:0]           axi_r_resp_o,
    output                  axi_r_user_o,
    output                  axi_r_last_o,
    output                  axi_r_valid_o,
    input                   axi_r_ready_i,

    // Regbus Request Input
    input wire [47:0]      reg_addr_i,
    input wire             reg_write_i,
    input wire [31:0]      reg_wdata_i,
    input wire [5:0]       reg_wstrb_i,
    input wire             reg_valid_i,

    // Regbus Request Output
    output wire            reg_error_o,
    output wire [31:0]     reg_rdata_o,
    output wire            reg_ready_o,

    // Controller to RPC DRAM Port
    output wire rpc_clk_o,
    output wire rpc_clk_no,
    output wire rpc_cs_no,
    output wire rpc_stb_o,

    inout  wire rpc_dqs,
    inout  wire rpc_dqsn,
    inout  wire rpc_db0,
    inout  wire rpc_db1,
    inout  wire rpc_db2,
    inout  wire rpc_db3,
    inout  wire rpc_db4,
    inout  wire rpc_db5,
    inout  wire rpc_db6,
    inout  wire rpc_db7,
    inout  wire rpc_db8,
    inout  wire rpc_db9,
    inout  wire rpc_dba,
    inout  wire rpc_dbb,
    inout  wire rpc_dbc,
    inout  wire rpc_dbd,
    inout  wire rpc_dbe,
    inout  wire rpc_dbf
);

  rpc_fpga_top i_rpc_wrap (

    // common signals
    .clkp_i                  (clkp_i),
    .clkn_i                  (clkn_i),
    .rst_ni                  (rst_ni),

    // axi slave port
    .axi_aw_id_i             (axi_aw_id_i),
    .axi_aw_addr_i           (axi_aw_addr_i),
    .axi_aw_len_i            (axi_aw_len_i),
    .axi_aw_size_i           (axi_aw_size_i),
    .axi_aw_burst_i          (axi_aw_burst_i),
    .axi_aw_lock_i           (axi_aw_lock_i),
    .axi_aw_cache_i          (axi_aw_cache_i),
    .axi_aw_prot_i           (axi_aw_prot_i),
    .axi_aw_qos_i            (axi_aw_qos_i),
    .axi_aw_region_i         (axi_aw_region_i),
    .axi_aw_atop_i           (axi_aw_atop_i),
    .axi_aw_user_i           (axi_aw_user_i),
    .axi_aw_valid_i          (axi_aw_valid_i),
    .axi_aw_ready_o          (axi_aw_ready_o),
    .axi_w_data_i            (axi_w_data_i),
    .axi_w_strb_i            (axi_w_strb_i),
    .axi_w_last_i            (axi_w_last_i),
    .axi_w_user_i            (axi_w_user_i),
    .axi_w_valid_i           (axi_w_valid_i),
    .axi_w_ready_o           (axi_w_ready_o),
    .axi_b_id_o              (axi_b_id_o),
    .axi_b_resp_o            (axi_b_resp_o),
    .axi_b_user_o            (axi_b_user_o),
    .axi_b_valid_o           (axi_b_valid_o),
    .axi_b_ready_i           (axi_b_ready_i),
    .axi_ar_id_i             (axi_ar_id_i),
    .axi_ar_addr_i           (axi_ar_addr_i),
    .axi_ar_len_i            (axi_ar_len_i),
    .axi_ar_size_i           (axi_ar_size_i),
    .axi_ar_burst_i          (axi_ar_burst_i),
    .axi_ar_lock_i           (axi_ar_lock_i),
    .axi_ar_cache_i          (axi_ar_cache_i),
    .axi_ar_prot_i           (axi_ar_prot_i),
    .axi_ar_qos_i            (axi_ar_qos_i),
    .axi_ar_region_i         (axi_ar_region_i),
    .axi_ar_user_i           (axi_ar_user_i),
    .axi_ar_valid_i          (axi_ar_valid_i),
    .axi_ar_ready_o          (axi_ar_ready_o),
    .axi_r_id_o              (axi_r_id_o),
    .axi_r_data_o            (axi_r_data_o),
    .axi_r_resp_o            (axi_r_resp_o),
    .axi_r_last_o            (axi_r_last_o),
    .axi_r_user_o            (axi_r_user_o),
    .axi_r_valid_o           (axi_r_valid_o),
    .axi_r_ready_i           (axi_r_ready_i),

    // Regbus Request Input
    .reg_addr_i              (reg_addr_i),
    .reg_write_i             (reg_write_i),
    .reg_wdata_i             (reg_wdata_i),
    .reg_wstrb_i             (reg_wstrb_i),
    .reg_valid_i             (reg_valid_i),

    // Regbus Request Output
    .reg_error_o             (reg_error_o),
    .reg_rdata_o             (reg_rdata_o),
    .reg_ready_o             (reg_ready_o),

    // Controller to RPC DRAM Port
    .rpc_clk_o               (rpc_clk_o),
    .rpc_clk_no              (rpc_clk_no),
    .rpc_cs_no               (rpc_cs_no),
    .rpc_stb_o               (rpc_stb_o),
    .rpc_dqs                 (rpc_dqs),
    .rpc_dqsn                (rpc_dqsn),
    .rpc_db0                 (rpc_db0),
    .rpc_db1                 (rpc_db1),
    .rpc_db2                 (rpc_db2),
    .rpc_db3                 (rpc_db3),
    .rpc_db4                 (rpc_db4),
    .rpc_db5                 (rpc_db5),
    .rpc_db6                 (rpc_db6),
    .rpc_db7                 (rpc_db7),
    .rpc_db8                 (rpc_db8),
    .rpc_db9                 (rpc_db9),
    .rpc_dba                 (rpc_dba),
    .rpc_dbb                 (rpc_dbb),
    .rpc_dbc                 (rpc_dbc),
    .rpc_dbd                 (rpc_dbd),
    .rpc_dbe                 (rpc_dbe),
    .rpc_dbf                 (rpc_dbf)
  );

endmodule
